module mdff(mout, min, mclk, mrst);

  input min, mclk, mrst;
  output mout;
  wire min, mclk, mrst;
  reg mout;
  
endmodule
